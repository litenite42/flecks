module main

import ecs
import util as u
//import ecs.managers as mgrs

fn main() {
	println('hello')

	mut coord := ecs.Coordinator{}
	dump(coord)
}
