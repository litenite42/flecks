module ecs