module ecs

import bitfield as bf

pub type Entity = i16
pub type ComponentType = i8

pub type Signature = bf.BitField
