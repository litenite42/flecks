module ecs

pub const (
	max_components = 32
	max_entities   = 5000
)
