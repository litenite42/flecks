module ecs
